library ieee;
use ieee.std_logic_1164.all;


entity latch_sre_nand is

	port (
	    S : in std_logic;
	    R : in std_logic;

        E : in std_logic;

        Q  : out std_logic;
        NQ : out std_logic
	    );

end entity;


architecture behavior of latch_sre_nand is

signal T  : std_logic;
signal NT : std_logic;

begin

    T  <= (S nand E) nand NT;
    NT <= (R nand E) nand T;

    Q  <= T;
    NQ <= NT;

end architecture;
